----------------------------------------------------------------------------------
--------------Visualizar Los Numeros En EL 7 Segmentos----------------------------
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity dis is
    Port ( Num1  : in  STD_LOGIC;
           Num2  : in  STD_LOGIC;
           Num3  : in  STD_LOGIC;
           Out1  : out STD_LOGIC;
           Out2  : out STD_LOGIC;
           Out3  : out STD_LOGIC;
           CLOCK : in  STD_LOGIC;
           RESET : in  STD_LOGIC);
end dis;

architecture Behavioral of dis is



begin


end Behavioral;

